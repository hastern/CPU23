library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;

entity E_ALU_ONEHOT is

    port (
        inp : in OpCode23;

        res : out Word23
    );

end entity;

architecture A_ALU_ONEHOT of E_ALU_ONEHOT is

begin
    process (inp)
    begin
        case inp is
            when "00000" => res <= "000000000000000000000000";
            when "00001" => res <= "000000000000000000000001";
            when "00010" => res <= "000000000000000000000010";
            when "00011" => res <= "000000000000000000000100";
            when "00100" => res <= "000000000000000000001000";
            when "00101" => res <= "000000000000000000010000";
            when "00110" => res <= "000000000000000000100000";
            when "00111" => res <= "000000000000000001000000";
            when "01000" => res <= "000000000000000010000000";
            when "01001" => res <= "000000000000000100000000";
            when "01010" => res <= "000000000000001000000000";
            when "01011" => res <= "000000000000010000000000";
            when "01100" => res <= "000000000000100000000000";
            when "01101" => res <= "000000000001000000000000";
            when "01110" => res <= "000000000010000000000000";
            when "01111" => res <= "000000000100000000000000";
            when "10000" => res <= "000000001000000000000000";
            when "10001" => res <= "000000010000000000000000";
            when "10010" => res <= "000000100000000000000000";
            when "10011" => res <= "000001000000000000000000";
            when "10100" => res <= "000010000000000000000000";
            when "10101" => res <= "000100000000000000000000";
            when "10110" => res <= "001000000000000000000000";
            when "10111" => res <= "010000000000000000000000";
            when "11000" => res <= "100000000000000000000000";
            when others  => res <= "000000000000000000000000";
        end case;
    end process;
end;
